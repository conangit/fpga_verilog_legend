module reverse_bits (
    input [7:0] a,
    output [0:7] b
    );
    
    assign b = a;
    
endmodule
